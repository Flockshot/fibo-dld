library verilog;
use verilog.vl_types.all;
entity Decoder_2_To_4_vlg_vec_tst is
end Decoder_2_To_4_vlg_vec_tst;
