module Dflip_tb();
  reg   Clk;
  reg   [3:0]D;
  wire  [3:0] Q;
  
  Dflip DUT (Q,D,Clk);
  always
  begin
    Clk=1; #50; 
    Clk=0; #50;
  end
  initial 
  begin
    D=4'b0000; #100;
    D=4'b0010; #100;
    D=4'b0100; #100;
    D=4'b1101; #100;
  end
endmodule

