module mux4to1_tb();
  parameter   size = 4;
  reg         [size-1:0]I1,I2,I3,I4;
  reg         [1:0]S;
  wire        [size-1:0]Y;
  mux4to1 DUT(I1,I2,I3,I4,S,Y);
  initial 
  begin
    I1=4'b0100; I2=4'b0010; I3=4'b1111; I4=4'b0000; S=2'b00; #100;
    I1=4'b0100; I2=4'b1110; I3=4'b0111; I4=4'b0010; S=2'b01; #100;
    I1=4'b0101; I2=4'b0010; I3=4'b1011; I4=4'b1100; S=2'b10; #100;
    I1=4'b1100; I2=4'b1010; I3=4'b1101; I4=4'b1000; S=2'b11; #100;
    
  end
endmodule
  




