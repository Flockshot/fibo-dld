module FIBO_DATAPATH_N (wrt_addr,wrt_en,clk,load_data,rd_addr1,rd_addr2,alu_opcode,count,zero_flag,data);
parameter size=4;
input wrt_en, clk, load_data;
input [1: 0] wrt_addr, rd_addr1, rd_addr2;
input [2: 0] alu_opcode;
input [size-1: 0] count;
output zero_flag;
output  [size-1: 0] data;
wire [3: 0] w1,w2;
wire [size-1:0] w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14;
decoder A1(wrt_addr, w1);
and (w2[3], w1[3], wrt_en);
and (w2[2], w1[2], wrt_en);
and (w2[1], w1[1], wrt_en);
and (w2[0], w1[0], wrt_en);
mux C1(data,count,load_data,w3); 
mux U0(w8,w3,w2[0],w4); 
mux U1(w9,w3,w2[1],w5);
mux U2(w10,w3,w2[2],w6);
mux U3(w11,w3,w2[3],w7);
Dflip D0(w8, w4, clk);
Dflip D1(w9, w5, clk);
Dflip D2(w10, w6, clk);
Dflip D3(w11, w7, clk);
mux4to1 B1(w8,w9,w10,w11,rd_addr1,w12); 
mux4to1 B2(w8,w9,w10,w11,rd_addr2,w13);  
ALU M1(w12,w13,alu_opcode,data,zero_flag);
Dflip D4(data,w14,clk);
endmodule
