library verilog;
use verilog.vl_types.all;
entity D_Flip_Flop_vlg_vec_tst is
end D_Flip_Flop_vlg_vec_tst;
