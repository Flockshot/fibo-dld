library verilog;
use verilog.vl_types.all;
entity Dflip_tb is
end Dflip_tb;
