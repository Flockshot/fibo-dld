library verilog;
use verilog.vl_types.all;
entity Four_Bit_4_To_1_Mux_vlg_vec_tst is
end Four_Bit_4_To_1_Mux_vlg_vec_tst;
