module Fibo_datapath_tb1();
parameter size=4;
reg wrt_en, clk, load_data;
reg [1:0] wrt_addr, rd_addr1, rd_addr2;
reg [2: 0] alu_opcode;
reg [size-1: 0] count;
wire zero_flag;
wire [size-1: 0] data;
FIBO_DATAPATH DUT(wrt_addr,wrt_en,clk,load_data,rd_addr1,rd_addr2,alu_opcode,count,zero_flag,data);
  always begin
  clk = 0; #25; clk = 1; #25; end
initial
 begin
   // R1 -> 01, R2 -> 10, R3-> 11, R4 = count -> 00
   //load count
  wrt_en=1;  load_data=1; wrt_addr=2'b00; rd_addr1=2'b00; rd_addr2=2'b00; alu_opcode=3'b100; count=4'b0110; #100;
  //set num1 and num2 (num1=num2=1)
  wrt_en=1;  load_data=0; wrt_addr=2'b01; rd_addr1=2'b01; rd_addr2=2'b01; alu_opcode=3'b001; count=4'b0110; #100;
  wrt_en=1;  load_data=0; wrt_addr=2'b10; rd_addr1=2'b10; rd_addr2=2'b10; alu_opcode=3'b001; count=4'b0110; #100;
  
  //R3<-R1
  wrt_en=1;  load_data=0; wrt_addr=2'b11; rd_addr1=2'b01; rd_addr2=2'b01; alu_opcode=3'b111; count=4'b0110; #100;
    //R1<-R1+R2
  wrt_en=1;  load_data=0; wrt_addr=2'b01; rd_addr1=2'b01; rd_addr2=2'b10; alu_opcode=3'b110; count=4'b0110; #100;
  //R2<-R3
  wrt_en=1;  load_data=0; wrt_addr=2'b10; rd_addr1=2'b11; rd_addr2=2'b11; alu_opcode=3'b111; count=4'b0110; #100;
  
   //R3<-R1
  wrt_en=1;  load_data=0; wrt_addr=2'b11; rd_addr1=2'b01; rd_addr2=2'b01; alu_opcode=3'b111; count=4'b0110; #100;
    //R1<-R1+R2
  wrt_en=1;  load_data=0; wrt_addr=2'b01; rd_addr1=2'b01; rd_addr2=2'b10; alu_opcode=3'b110; count=4'b0110; #100;
  //R2<-R3
  wrt_en=1;  load_data=0; wrt_addr=2'b10; rd_addr1=2'b11; rd_addr2=2'b11; alu_opcode=3'b111; count=4'b0110; #100;
  
  //R3<-R1
  wrt_en=1;  load_data=0; wrt_addr=2'b11; rd_addr1=2'b01; rd_addr2=2'b01; alu_opcode=3'b111; count=4'b0110; #100;
    //R1<-R1+R2
  wrt_en=1;  load_data=0; wrt_addr=2'b01; rd_addr1=2'b01; rd_addr2=2'b10; alu_opcode=3'b110; count=4'b0110; #100;
  //R2<-R3
  wrt_en=1;  load_data=0; wrt_addr=2'b10; rd_addr1=2'b11; rd_addr2=2'b11; alu_opcode=3'b111; count=4'b0110; #100;
  
  //R3<-R1
  wrt_en=1;  load_data=0; wrt_addr=2'b11; rd_addr1=2'b01; rd_addr2=2'b01; alu_opcode=3'b111; count=4'b0110; #100;
    //R1<-R1+R2
  wrt_en=1;  load_data=0; wrt_addr=2'b01; rd_addr1=2'b01; rd_addr2=2'b10; alu_opcode=3'b110; count=4'b0110; #100;
  //R2<-R3
  wrt_en=1;  load_data=0; wrt_addr=2'b10; rd_addr1=2'b11; rd_addr2=2'b11; alu_opcode=3'b111; count=4'b0110; #100;
  
//R3<-R1
  wrt_en=1;  load_data=0; wrt_addr=2'b11; rd_addr1=2'b01; rd_addr2=2'b01; alu_opcode=3'b111; count=4'b0110; #100;
    //R1<-R1+R2
  wrt_en=1;  load_data=0; wrt_addr=2'b01; rd_addr1=2'b01; rd_addr2=2'b10; alu_opcode=3'b110; count=4'b0110; #100;
  //R2<-R3
  wrt_en=1;  load_data=0; wrt_addr=2'b10; rd_addr1=2'b11; rd_addr2=2'b11; alu_opcode=3'b111; count=4'b0110; #100;
  end
  endmodule

